interface gpio_if;

  logic clk;
  logic[31:0] gpio;
  bit ext_clk;

endinterface: gpio_if
